library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity floppy_burt_top is
    port (
        CLOCK_50 : in std_logic;
        VGA_R, VGA_G, VGA_B : out std_logic_vector(3 downto 0);
        VGA_HS, VGA_VS : out std_logic
    );
end floppy_burt_top; 

architecture vga_test of floppy_burt_top is

    component VGA_SYNC is
        port (
            clock_25Mhz : in STD_LOGIC; 
            red, green, blue : in STD_LOGIC_VECTOR(3 downto 0);
            red_out, green_out, blue_out : out STD_LOGIC_VECTOR(3 downto 0);
            horiz_sync_out, vert_sync_out : out STD_LOGIC;
            pixel_row, pixel_column: out STD_LOGIC_VECTOR(9 downto 0)
        );
    end component VGA_SYNC;

    component ball IS
        port (
            clk : in std_logic;
            pixel_row, pixel_column	: in std_logic_vector(9 downto 0);
            red, green, blue : out std_logic_vector(3 downto 0)
        );		
    end component ball;

    component pll25MHz is
        port (
            refclk   : in  std_logic := '0'; --  refclk.clk
            rst      : in  std_logic := '0'; --   reset.reset
            outclk_0 : out std_logic;        -- outclk0.clk
            locked   : out std_logic         --  locked.export
        );
    end component pll25MHz;

    -- INTERMEDIATE SIGNALS
    signal clock_25Mhz : std_logic;
    signal s_rst : std_logic; -- can link to board reset if want
    signal s_locked : std_logic; -- ? clock stability

    signal s_pix_row : std_logic_vector(9 downto 0);
    signal s_pix_col : std_logic_vector(9 downto 0);
    signal s_red : std_logic_vector(3 downto 0);
    signal s_green : std_logic_vector(3 downto 0);
    signal s_blue : std_logic_vector(3 downto 0);

    -- need to know fpga pin ports:
    -- for sync and colors

begin

c1: pll25MHz
    port map (
        refclk => CLOCK_50,
        rst => s_rst,
        outclk_0 => clock_25Mhz,
        locked => s_locked
    );

b1: ball
    port map (
        -- input
        clk => clock_25Mhz,
        pixel_row => s_pix_row,
        pixel_column => s_pix_col,
        -- output
        red => s_red,
        green => s_green,
        blue => s_blue
    );

v1: VGA_SYNC
    port map (
        -- input
        clock_25Mhz => clock_25Mhz,
        red => s_red,
        green => s_green,
        blue => s_blue,
        -- output
        -- NOTE: might have to do a different approach for the color mapping - but just test it first
        -- if not working then just make it the entire stdlogicvector, but check ball to see if changes needed
        red_out => VGA_R, 
        green_out => VGA_G,
        blue_out => VGA_B,
        horiz_sync_out => VGA_HS,
        vert_sync_out => VGA_VS,
        pixel_row => s_pix_row, 
        pixel_column => s_pix_col
    );

end architecture;